module	Lab_0	(a,b,c);

input a,b;
output c;

assign	c	=	a&b;

endmodule

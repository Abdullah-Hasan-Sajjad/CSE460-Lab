module	exp2(w,,presentState,nextState,clock,reset);

endmodule
module	Lab2_assessment(w,y)

input [3:0]w;
output reg[1:0]y;



endmodule